library verilog;
use verilog.vl_types.all;
entity receive_top_module_tb is
end receive_top_module_tb;
