library verilog;
use verilog.vl_types.all;
entity butterfly_radix4_2nd is
    generic(
        cos0            : integer := 32767;
        cos1            : integer := 32767;
        cos2            : integer := 32767;
        cos3            : integer := 30273;
        cos4            : integer := 23170;
        cos5            : integer := 12540;
        cos6            : integer := 23170;
        cos7            : integer := 0;
        cos8            : integer := 42366;
        cos9            : integer := 12540;
        cos10           : integer := 42366;
        cos11           : integer := 35263;
        sin0            : integer := 0;
        sin1            : integer := 0;
        sin2            : integer := 0;
        sin3            : integer := 52996;
        sin4            : integer := 42366;
        sin5            : integer := 35263;
        sin6            : integer := 42366;
        sin7            : integer := 32769;
        sin8            : integer := 42366;
        sin9            : integer := 35263;
        sin10           : integer := 42366;
        sin11           : integer := 12540
    );
    port(
        clk             : in     vl_logic;
        re_0            : in     vl_logic_vector(15 downto 0);
        re_1            : in     vl_logic_vector(15 downto 0);
        re_2            : in     vl_logic_vector(15 downto 0);
        re_3            : in     vl_logic_vector(15 downto 0);
        re_4            : in     vl_logic_vector(15 downto 0);
        re_5            : in     vl_logic_vector(15 downto 0);
        re_6            : in     vl_logic_vector(15 downto 0);
        re_7            : in     vl_logic_vector(15 downto 0);
        re_8            : in     vl_logic_vector(15 downto 0);
        re_9            : in     vl_logic_vector(15 downto 0);
        re_10           : in     vl_logic_vector(15 downto 0);
        re_11           : in     vl_logic_vector(15 downto 0);
        re_12           : in     vl_logic_vector(15 downto 0);
        re_13           : in     vl_logic_vector(15 downto 0);
        re_14           : in     vl_logic_vector(15 downto 0);
        re_15           : in     vl_logic_vector(15 downto 0);
        im_0            : in     vl_logic_vector(15 downto 0);
        im_1            : in     vl_logic_vector(15 downto 0);
        im_2            : in     vl_logic_vector(15 downto 0);
        im_3            : in     vl_logic_vector(15 downto 0);
        im_4            : in     vl_logic_vector(15 downto 0);
        im_5            : in     vl_logic_vector(15 downto 0);
        im_6            : in     vl_logic_vector(15 downto 0);
        im_7            : in     vl_logic_vector(15 downto 0);
        im_8            : in     vl_logic_vector(15 downto 0);
        im_9            : in     vl_logic_vector(15 downto 0);
        im_10           : in     vl_logic_vector(15 downto 0);
        im_11           : in     vl_logic_vector(15 downto 0);
        im_12           : in     vl_logic_vector(15 downto 0);
        im_13           : in     vl_logic_vector(15 downto 0);
        im_14           : in     vl_logic_vector(15 downto 0);
        im_15           : in     vl_logic_vector(15 downto 0);
        butterfly_re0   : out    vl_logic_vector(15 downto 0);
        butterfly_re1   : out    vl_logic_vector(15 downto 0);
        butterfly_re2   : out    vl_logic_vector(15 downto 0);
        butterfly_re3   : out    vl_logic_vector(15 downto 0);
        butterfly_re4   : out    vl_logic_vector(15 downto 0);
        butterfly_re5   : out    vl_logic_vector(15 downto 0);
        butterfly_re6   : out    vl_logic_vector(15 downto 0);
        butterfly_re7   : out    vl_logic_vector(15 downto 0);
        butterfly_re8   : out    vl_logic_vector(15 downto 0);
        butterfly_re9   : out    vl_logic_vector(15 downto 0);
        butterfly_re10  : out    vl_logic_vector(15 downto 0);
        butterfly_re11  : out    vl_logic_vector(15 downto 0);
        butterfly_re12  : out    vl_logic_vector(15 downto 0);
        butterfly_re13  : out    vl_logic_vector(15 downto 0);
        butterfly_re14  : out    vl_logic_vector(15 downto 0);
        butterfly_re15  : out    vl_logic_vector(15 downto 0);
        butterfly_im0   : out    vl_logic_vector(15 downto 0);
        butterfly_im1   : out    vl_logic_vector(15 downto 0);
        butterfly_im2   : out    vl_logic_vector(15 downto 0);
        butterfly_im3   : out    vl_logic_vector(15 downto 0);
        butterfly_im4   : out    vl_logic_vector(15 downto 0);
        butterfly_im5   : out    vl_logic_vector(15 downto 0);
        butterfly_im6   : out    vl_logic_vector(15 downto 0);
        butterfly_im7   : out    vl_logic_vector(15 downto 0);
        butterfly_im8   : out    vl_logic_vector(15 downto 0);
        butterfly_im9   : out    vl_logic_vector(15 downto 0);
        butterfly_im10  : out    vl_logic_vector(15 downto 0);
        butterfly_im11  : out    vl_logic_vector(15 downto 0);
        butterfly_im12  : out    vl_logic_vector(15 downto 0);
        butterfly_im13  : out    vl_logic_vector(15 downto 0);
        butterfly_im14  : out    vl_logic_vector(15 downto 0);
        butterfly_im15  : out    vl_logic_vector(15 downto 0)
    );
end butterfly_radix4_2nd;
