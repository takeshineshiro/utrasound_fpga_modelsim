
  

 module  cc3200_model_gen   (
 //input
    input         clk_in ,
    input         reset_n
//output
     

 );







 endmodule 
  
