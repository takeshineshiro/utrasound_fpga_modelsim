
module   cmd_gen_submodule (



);




endmodule
