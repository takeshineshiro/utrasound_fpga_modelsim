
  module   data_gen_submodule  (
     //input
           input                  clk     ,

           input                  reset_n , 
              
      //output
          output  [11:0]          Data_A  ,

          output  [11:0]          Data_B  ,

          output  [11:0]          Data_C  ,

          output  [11:0]          Data_D  ,
              
          output  [11:0]          Data_E  ,

          output  [11:0]          Data_F  ,  
       
          output  [11:0]          Data_G  ,

          output  [11:0]          Data_H     
              


  );











endmodule
