library verilog;
use verilog.vl_types.all;
entity transmit_test_entity_tb is
end transmit_test_entity_tb;
